.TITLE FUZZ - FREQUENCY RESPONSE

.INCLUDE 1N4148_DI.model
.INCLUDE BC107.model

VCC 5 0 9
VCC 7 0 9

V1 1 0 DC 0 AC 1

C1 3 4 50n
C2 6 8 1500p
C3 8 9 50n

R1 1 2 470k
R2a 2 3 1K
R2b 3 0 99k
R3 4 6 2200k
R4 5 6 100k
R5 6 8 2200k
R6 7 8 100k
R7 9 0 100k

D1 9 0 1N4148_DI
D2 0 9 1N4148_DI

Q1 6 4 0 BC107
Q2 8 6 0 BC107


.PRINT OP Iter(0) V(3)

.PRINT AC VDB(9)

*     FROM      TO   STEP
.TRAN 0.00001   0.2  0.0001

*       #STEPS/DECADE FROM   TO 
.AC DEC 20            0.1    10Meg

.END
